library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package program is
    type program_t is array(0 to 1023) of unsigned(31 downto 0);

    constant program_c: program_t := (

        -- 0: movhi r1, b"0000000000010000"
        b"000100_00001_0000000000010000_00000",

        -- 1: subi r1, r1, 1
        b"001101_00001_00001_0000000000000001",

        -- 2: cmpi r1, 0
        b"100100_00000_00001_0000000000000000",

        -- 3: bneq -3
        b"101001_11111111111111111111111101",

        -- 4: addi r2, r0, b"0000000011111111"
        b"001011_00010_00000_0000000011111111",

        -- 5: str r0, r2, 1024
        b"000010_00000_00000_00010_10000000000",

        -- 6: movhi r1, b"0000000000010000"
        b"000100_00001_0000000000010000_00000",

        -- 7: subi r1, r1, 1
        b"001101_00001_00001_0000000000000001",

        -- 8: cmpi r1, 0
        b"100100_00000_00001_0000000000000000",

        -- 9: bneq -3
        b"101001_11111111111111111111111101",

        -- 10: add r2, r0, r0
        b"001010_00010_00000_00000_00000000000",

        -- 11: str r0, r2, 1024
        b"000010_00000_00000_00010_10000000000",

        -- 12: jmp r0, 0
        b"101110_00000_00000_0000000000000000",

        others => (others => '0')
    );
end program;
